module xor_gate(input wire [19:0] a, input wire [19:0] b, output wire [19:0] c);

    assign c = a^b;

endmodule