module not_gate(input wire [19:0] a, output wire [19:0] b);

    assign b = ~a;

endmodule