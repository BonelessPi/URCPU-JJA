module increment_module(input wire [19:0] in, output wire [19:0] out);

    assign out = in+1;

endmodule